--writeToSDComponent